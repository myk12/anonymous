`resetall
`timescale 1ns / 1ps
`default_nettype none

/*
 * Time synchronization master module
 */
module time_sync_master #
(
    parameter SYNC_TS_WIDTH = 32,
    parameter IDENTIFIER_WIDTH = 16,
    parameter PORT_ID_WIDTH = 4,

    // self ID
    parameter SELF_ID = 123456,

    // AXIS interface
    parameter AXIS_DATA_WIDTH = 64,
    parameter AXIS_KEEP_WIDTH = (AXIS_DATA_WIDTH/8),
    parameter AXIS_TX_ID_WIDTH = 8,
    parameter AXIS_TX_DEST_WIDTH = 8,
    parameter AXIS_TX_USER_WIDTH = 1
)
(
    input wire                                      clk,
    input wire                                      rst,

    // time stamp input
    input wire [95:0]                               ptp_ts_tod,

    // sync scheduler output
    input wire                                      sync_enable,
    input wire [IDENTIFIER_WIDTH-1:0]               sync_dest_id,

    // master sync packet output
    output wire [AXIS_DATA_WIDTH-1:0]               m_axis_sync_tx_data,
    output wire [AXIS_KEEP_WIDTH-1:0]               m_axis_sync_tx_keep,
    output wire                                     m_axis_sync_tx_valid,
    input wire                                      m_axis_sync_tx_ready,
    output wire                                     m_axis_sync_tx_last,
    output wire [AXIS_TX_ID_WIDTH-1:0]              m_axis_sync_tx_id,
    output wire [AXIS_TX_DEST_WIDTH-1:0]            m_axis_sync_tx_dest,
    output wire [AXIS_TX_USER_WIDTH-1:0]            m_axis_sync_tx_user,

    // time sync TX checksum command
    output wire                                     sync_tx_csum_cmd_csum_enable,
    output wire [7:0]                               sync_tx_csum_cmd_csum_start,
    output wire [7:0]                               sync_tx_csum_cmd_csum_offset,
    output wire                                     sync_tx_csum_cmd_valid,
    input wire                                      sync_tx_csum_cmd_ready 
);
//
// Info: This module is a time synchronization master module that sends time synchronization packets
// to the time synchronization slave module. It receives the timestamp from the PTP and is enabled
// by the sync_enable signal that is generated by the time synchronization scheduler module.

// define the state machine
parameter STATE_IDLE        = 0;
parameter STATE_CSUM_ENABLE = 1;
parameter STATE_WAIT_READY  = 2;
parameter STATE_TX_DATA     = 3;

reg [1:0] state, next_state;

reg sync_enable_reg;
reg [IDENTIFIER_WIDTH-1:0] sync_dest_reg;

// AXI stream signals
reg [AXIS_DATA_WIDTH-1:0]       tx_data_reg;
reg [AXIS_KEEP_WIDTH-1:0]       tx_keep_reg;
reg                             tx_valid_reg;
reg                             tx_last_reg;
reg [AXIS_TX_ID_WIDTH-1:0]      tx_id_reg;
reg [AXIS_TX_DEST_WIDTH-1:0]    tx_dest_reg;
reg [AXIS_TX_USER_WIDTH-1:0]    tx_user_reg;

// TX checksum command
reg             tx_csum_cmd_csum_enable_reg;
reg [7:0]       tx_csum_cmd_csum_start_reg;
reg [7:0]       tx_csum_cmd_csum_offset_reg;
reg             tx_csum_cmd_valid_reg;

assign m_axis_sync_tx_data  = tx_data_reg;
assign m_axis_sync_tx_keep  = tx_keep_reg;
assign m_axis_sync_tx_valid = tx_valid_reg;
assign m_axis_sync_tx_last  = tx_last_reg;
assign m_axis_sync_tx_id    = tx_id_reg;
assign m_axis_sync_tx_dest  = tx_dest_reg;
assign m_axis_sync_tx_user  = tx_user_reg;

assign sync_tx_csum_cmd_csum_enable = tx_csum_cmd_csum_enable_reg;
assign sync_tx_csum_cmd_csum_start  = tx_csum_cmd_csum_start_reg;
assign sync_tx_csum_cmd_csum_offset = tx_csum_cmd_csum_offset_reg;
assign sync_tx_csum_cmd_valid       = tx_csum_cmd_valid_reg;

// state machine
always @(*) begin
    case (state)
        STATE_IDLE : begin
            if (sync_enable_reg) begin
                next_state = STATE_CSUM_ENABLE;
            end else begin
                next_state = STATE_IDLE;
            end
        end
        STATE_CSUM_ENABLE: begin
            next_state = STATE_WAIT_READY;
        end
        STATE_WAIT_READY: begin
            if (m_axis_sync_tx_ready) begin
                next_state = STATE_TX_DATA;
            end else begin
                next_state = STATE_WAIT_READY;
            end
        end
        STATE_TX_DATA: begin
            next_state = STATE_IDLE;
        end
        default: next_state = STATE_IDLE;
    endcase
end

// state transition
always @(posedge clk or posedge rst) begin
    if (rst) begin
        state <= STATE_IDLE;
    end else begin
        state <= next_state;
    end
end

always @(posedge clk or posedge rst) begin
    if (rst) begin
        sync_enable_reg <= 0;
        sync_dest_reg <= 0;

        tx_data_reg <= 0;
        tx_keep_reg <= 0;
        tx_valid_reg <= 0;
        tx_last_reg <= 0;
        tx_id_reg <= 0;
        tx_dest_reg <= 0;
        tx_user_reg <= 0;
        tx_csum_cmd_csum_enable_reg <= 0;
        tx_csum_cmd_csum_start_reg <= 0;
        tx_csum_cmd_csum_offset_reg <= 0;
        tx_csum_cmd_valid_reg <= 0;
    end else begin
        case (state)
            STATE_IDLE: begin
                sync_enable_reg <= sync_enable;
                sync_dest_reg <= sync_dest_id;

                tx_data_reg <= 0;
                tx_keep_reg <= 0;
                tx_valid_reg <= 0;
                tx_last_reg <= 0;
                tx_id_reg <= 0;
                tx_dest_reg <= 0;
                tx_user_reg <= 0;

                tx_csum_cmd_csum_enable_reg <= 0;
                tx_csum_cmd_csum_start_reg <= 0;
                tx_csum_cmd_csum_offset_reg <= 0;
                tx_csum_cmd_valid_reg <= 0;
            end
            STATE_CSUM_ENABLE: begin
                sync_enable_reg <= 0;

                tx_csum_cmd_csum_enable_reg <= 0;
                tx_csum_cmd_csum_start_reg <= 0;
                tx_csum_cmd_csum_offset_reg <= 0;
                tx_csum_cmd_valid_reg <= 1;
            end
            STATE_WAIT_READY: begin
                // Generate the sync packet
                // format:
                // [15:0] magic: 0x77f8
                // [31:16] dest: sync_dest_reg
                // [47:32] src:  0x1176
                // [143:48] timestamp: ptp_ts_tod[95:0]
                tx_data_reg[15:0] <= 16'h77f8;
                tx_data_reg[31:16] <= sync_dest_reg;
                tx_data_reg[47:32] <= 16'h1176;
                tx_data_reg[143:48] <= ptp_ts_tod;
                tx_keep_reg <= {AXIS_KEEP_WIDTH{1'b1}};
                tx_id_reg <= 1;
                tx_dest_reg <= 1;
                tx_user_reg <= 0;

                tx_csum_cmd_csum_enable_reg <= 0;
                tx_csum_cmd_csum_start_reg <= 0;
                tx_csum_cmd_csum_offset_reg <= 0;
                tx_csum_cmd_valid_reg <= 0;
            end
            STATE_TX_DATA: begin
                tx_data_reg <= tx_data_reg;
                tx_keep_reg <= tx_keep_reg;
                tx_valid_reg <= 1;
                tx_last_reg <= 1;
                tx_id_reg <= tx_id_reg;
                tx_dest_reg <= tx_dest_reg;
                tx_user_reg <= tx_user_reg;

                tx_csum_cmd_csum_enable_reg <= 0;
                tx_csum_cmd_csum_start_reg <= 0;
                tx_csum_cmd_csum_offset_reg <= 0;
                tx_csum_cmd_valid_reg <= 0;
            end
            default: begin
                sync_enable_reg <= 0;
                tx_data_reg <= 0;
                tx_keep_reg <= 0;
                tx_valid_reg <= 0;
                tx_last_reg <= 0;
                tx_id_reg <= 0;
                tx_dest_reg <= 0;
                tx_user_reg <= 0;
                tx_csum_cmd_csum_enable_reg <= 0;
                tx_csum_cmd_csum_start_reg <= 0;
                tx_csum_cmd_csum_offset_reg <= 0;
                tx_csum_cmd_valid_reg <= 0;
            end
        endcase
    end
end

endmodule
